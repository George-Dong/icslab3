`ifndef __CPUHEAD_SVH__
`define __CPUHEAD_SVH__

`include "common.svh"
`include "cp0.svh"
`include "content.svh"

`endif
