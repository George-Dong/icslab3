`ifndef __REFCPU_DEFS_SVH__
`define __REFCPU_DEFS_SVH__

`include "common.svh"
`include "shortcut.svh"

`include "instr.svh"
`include "cp0.svh"
`include "context.svh"

`endif
